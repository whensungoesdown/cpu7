module mul32x32(
    input  wire [32:0] a,
    input  wire [32:0] b,
    input  wire        a_sign,
    input  wire        b_sign,
    output      [65:0] u,
    output      [65:0] v
);
wire [15:0] enc_ext  ;                        
wire        enc_lastb;                        
wire [16:0] enc_m1   ;                        
wire [16:0] enc_m2   ;                        
wire [16:0] enc_neg  ;                        
wire [65:0] tree_c0  ;                        
wire [65:0] tree_c1  ;                        
wire [65:0] tree_c10 ;                        
wire [65:0] tree_c11 ;                        
wire [65:0] tree_c12 ;                        
wire [65:0] tree_c13 ;                        
wire [65:0] tree_c14 ;                        
wire [65:0] tree_c15 ;                        
wire [65:0] tree_c2  ;                        
wire [65:0] tree_c3  ;                        
wire [65:0] tree_c4  ;                        
wire [65:0] tree_c5  ;                        
wire [65:0] tree_c6  ;                        
wire [65:0] tree_c7  ;                        
wire [65:0] tree_c8  ;                        
wire [65:0] tree_c9  ;                        
wire [65:0] tree_s0  ;                        
wire [65:0] tree_s1  ;                        
wire [65:0] tree_s10 ;                        
wire [65:0] tree_s11 ;                        
wire [65:0] tree_s12 ;                        
wire [65:0] tree_s13 ;                        
wire [65:0] tree_s14 ;                        
wire [65:0] tree_s15 ;                        
wire [65:0] tree_s2  ;                        
wire [65:0] tree_s3  ;                        
wire [65:0] tree_s4  ;                        
wire [65:0] tree_s5  ;                        
wire [65:0] tree_s6  ;                        
wire [65:0] tree_s7  ;                        
wire [65:0] tree_s8  ;                        
wire [65:0] tree_s9  ;                        
wire [32:0] y0       ;                        
wire [32:0] y1       ;                        
wire [32:0] y10      ;                        
wire [32:0] y11      ;                        
wire [32:0] y12      ;                        
wire [32:0] y13      ;                        
wire [32:0] y14      ;                        
wire [32:0] y15      ;                        
wire [32:0] y16      ;                        
wire [32:0] y2       ;                        
wire [32:0] y3       ;                        
wire [32:0] y4       ;                        
wire [32:0] y5       ;                        
wire [32:0] y6       ;                        
wire [32:0] y7       ;                        
wire [32:0] y8       ;                        
wire [32:0] y9       ;                        
wire [65:0] z0       ;                        
wire [65:0] z1       ;                        
wire [65:0] z10      ;                        
wire [65:0] z11      ;                        
wire [65:0] z12      ;                        
wire [65:0] z13      ;                        
wire [65:0] z14      ;                        
wire [65:0] z15      ;                        
wire [65:0] z16      ;                        
wire [65:0] z17      ;
wire [65:0] z2       ;                        
wire [65:0] z3       ;                        
wire [65:0] z4       ;                        
wire [65:0] z5       ;                        
wire [65:0] z6       ;                        
wire [65:0] z7       ;                        
wire [65:0] z8       ;                        
wire [65:0] z9       ;                        
assign enc_ext  [0 ] = enc_lastb && a[0] && !a[1] || !enc_lastb && a[1];
assign enc_ext  [1 ] = (a[1 ] || a[2 ]) && !a[3 ] && enc_lastb || !(a[1 ] && a[2 ]) && a[3 ] && !enc_lastb;
assign enc_ext  [2 ] = (a[3 ] || a[4 ]) && !a[5 ] && enc_lastb || !(a[3 ] && a[4 ]) && a[5 ] && !enc_lastb;
assign enc_ext  [3 ] = (a[5 ] || a[6 ]) && !a[7 ] && enc_lastb || !(a[5 ] && a[6 ]) && a[7 ] && !enc_lastb;
assign enc_ext  [4 ] = (a[7 ] || a[8 ]) && !a[9 ] && enc_lastb || !(a[7 ] && a[8 ]) && a[9 ] && !enc_lastb;
assign enc_ext  [5 ] = (a[9 ] || a[10]) && !a[11] && enc_lastb || !(a[9 ] && a[10]) && a[11] && !enc_lastb;
assign enc_ext  [6 ] = (a[11] || a[12]) && !a[13] && enc_lastb || !(a[11] && a[12]) && a[13] && !enc_lastb;
assign enc_ext  [7 ] = (a[13] || a[14]) && !a[15] && enc_lastb || !(a[13] && a[14]) && a[15] && !enc_lastb;
assign enc_ext  [8 ] = (a[15] || a[16]) && !a[17] && enc_lastb || !(a[15] && a[16]) && a[17] && !enc_lastb;
assign enc_ext  [9 ] = (a[17] || a[18]) && !a[19] && enc_lastb || !(a[17] && a[18]) && a[19] && !enc_lastb;
assign enc_ext  [10] = (a[19] || a[20]) && !a[21] && enc_lastb || !(a[19] && a[20]) && a[21] && !enc_lastb;
assign enc_ext  [11] = (a[21] || a[22]) && !a[23] && enc_lastb || !(a[21] && a[22]) && a[23] && !enc_lastb;
assign enc_ext  [12] = (a[23] || a[24]) && !a[25] && enc_lastb || !(a[23] && a[24]) && a[25] && !enc_lastb;
assign enc_ext  [13] = (a[25] || a[26]) && !a[27] && enc_lastb || !(a[25] && a[26]) && a[27] && !enc_lastb;
assign enc_ext  [14] = (a[27] || a[28]) && !a[29] && enc_lastb || !(a[27] && a[28]) && a[29] && !enc_lastb;
assign enc_ext  [15] = (a[29] || a[30]) && !a[31] && enc_lastb || !(a[29] && a[30]) && a[31] && !enc_lastb;
assign enc_lastb     = b_sign && b[32];
assign enc_m1   [0 ] = a[0];
assign enc_m1   [1 ] = a[1 ] ^ a[2 ];
assign enc_m1   [2 ] = a[3 ] ^ a[4 ];
assign enc_m1   [3 ] = a[5 ] ^ a[6 ];
assign enc_m1   [4 ] = a[7 ] ^ a[8 ];
assign enc_m1   [5 ] = a[9 ] ^ a[10];
assign enc_m1   [6 ] = a[11] ^ a[12];
assign enc_m1   [7 ] = a[13] ^ a[14];
assign enc_m1   [8 ] = a[15] ^ a[16];
assign enc_m1   [9 ] = a[17] ^ a[18];
assign enc_m1   [10] = a[19] ^ a[20];
assign enc_m1   [11] = a[21] ^ a[22];
assign enc_m1   [12] = a[23] ^ a[24];
assign enc_m1   [13] = a[25] ^ a[26];
assign enc_m1   [14] = a[27] ^ a[28];
assign enc_m1   [15] = a[29] ^ a[30];
assign enc_m1   [16] = a[32] ^ a[31];
assign enc_m2   [0 ] = a[1] && !a[0];
assign enc_m2   [1 ] = a[1 ] && a[2 ] && !a[3 ] || !a[1 ] && !a[2 ] && a[3 ];
assign enc_m2   [2 ] = a[3 ] && a[4 ] && !a[5 ] || !a[3 ] && !a[4 ] && a[5 ];
assign enc_m2   [3 ] = a[5 ] && a[6 ] && !a[7 ] || !a[5 ] && !a[6 ] && a[7 ];
assign enc_m2   [4 ] = a[7 ] && a[8 ] && !a[9 ] || !a[7 ] && !a[8 ] && a[9 ];
assign enc_m2   [5 ] = a[9 ] && a[10] && !a[11] || !a[9 ] && !a[10] && a[11];
assign enc_m2   [6 ] = a[11] && a[12] && !a[13] || !a[11] && !a[12] && a[13];
assign enc_m2   [7 ] = a[13] && a[14] && !a[15] || !a[13] && !a[14] && a[15];
assign enc_m2   [8 ] = a[15] && a[16] && !a[17] || !a[15] && !a[16] && a[17];
assign enc_m2   [9 ] = a[17] && a[18] && !a[19] || !a[17] && !a[18] && a[19];
assign enc_m2   [10] = a[19] && a[20] && !a[21] || !a[19] && !a[20] && a[21];
assign enc_m2   [11] = a[21] && a[22] && !a[23] || !a[21] && !a[22] && a[23];
assign enc_m2   [12] = a[23] && a[24] && !a[25] || !a[23] && !a[24] && a[25];
assign enc_m2   [13] = a[25] && a[26] && !a[27] || !a[25] && !a[26] && a[27];
assign enc_m2   [14] = a[27] && a[28] && !a[29] || !a[27] && !a[28] && a[29];
assign enc_m2   [15] = a[29] && a[30] && !a[31] || !a[29] && !a[30] && a[31];
assign enc_m2   [16] = a[32] && a[31] && !a_sign;
assign enc_neg  [0 ] = a[1];
assign enc_neg  [1 ] = a[3 ] && !(a[1 ] && a[2 ]);
assign enc_neg  [2 ] = a[5 ] && !(a[3 ] && a[4 ]);
assign enc_neg  [3 ] = a[7 ] && !(a[5 ] && a[6 ]);
assign enc_neg  [4 ] = a[9 ] && !(a[7 ] && a[8 ]);
assign enc_neg  [5 ] = a[11] && !(a[9 ] && a[10]);
assign enc_neg  [6 ] = a[13] && !(a[11] && a[12]);
assign enc_neg  [7 ] = a[15] && !(a[13] && a[14]);
assign enc_neg  [8 ] = a[17] && !(a[15] && a[16]);
assign enc_neg  [9 ] = a[19] && !(a[17] && a[18]);
assign enc_neg  [10] = a[21] && !(a[19] && a[20]);
assign enc_neg  [11] = a[23] && !(a[21] && a[22]);
assign enc_neg  [12] = a[25] && !(a[23] && a[24]);
assign enc_neg  [13] = a[27] && !(a[25] && a[26]);
assign enc_neg  [14] = a[29] && !(a[27] && a[28]);
assign enc_neg  [15] = a[31] && !(a[29] && a[30]);
assign enc_neg  [16] = a[32] && !a[31] && a_sign;
assign tree_c0       = {z0      [64:0] & z1      [64:0] | z0      [64:0] & z2      [64:0] | z1      [64:0] & z2      [64:0],1'b0};
assign tree_c1       = {z3      [64:0] & z4      [64:0] | z3      [64:0] & z5      [64:0] | z4      [64:0] & z5      [64:0],1'b0};
assign tree_c10      = {tree_s6 [64:0] & tree_s7 [64:0] | tree_s6 [64:0] & tree_s8 [64:0] | tree_s7 [64:0] & tree_s8 [64:0],1'b0};
assign tree_c11      = {tree_s9 [64:0] & tree_c6 [64:0] | tree_s9 [64:0] & tree_c7 [64:0] | tree_c6 [64:0] & tree_c7 [64:0],1'b0};
assign tree_c12      = {tree_c8 [64:0] & tree_c9 [64:0] | tree_c8 [64:0] & tree_s10[64:0] | tree_c9 [64:0] & tree_s10[64:0],1'b0};
assign tree_c13      = {tree_s11[64:0] & tree_c10[64:0] | tree_s11[64:0] & tree_c11[64:0] | tree_c10[64:0] & tree_c11[64:0],1'b0};
assign tree_c14      = {tree_s12[64:0] & tree_s13[64:0] | tree_s12[64:0] & tree_c12[64:0] | tree_s13[64:0] & tree_c12[64:0],1'b0};
assign tree_c15      = {tree_c13[64:0] & tree_s14[64:0] | tree_c13[64:0] & tree_c14[64:0] | tree_s14[64:0] & tree_c14[64:0],1'b0};
assign tree_c2       = {z6      [64:0] & z7      [64:0] | z6      [64:0] & z8      [64:0] | z7      [64:0] & z8      [64:0],1'b0};
assign tree_c3       = {z9      [64:0] & z10     [64:0] | z9      [64:0] & z11     [64:0] | z10     [64:0] & z11     [64:0],1'b0};
assign tree_c4       = {z12     [64:0] & z13     [64:0] | z12     [64:0] & z14     [64:0] | z13     [64:0] & z14     [64:0],1'b0};
assign tree_c5       = {z15     [64:0] & z16     [64:0] | z15     [64:0] & z17     [64:0] | z16     [64:0] & z17     [64:0],1'b0};
assign tree_c6       = {tree_s0 [64:0] & tree_s1 [64:0] | tree_s0 [64:0] & tree_s2 [64:0] | tree_s1 [64:0] & tree_s2 [64:0],1'b0};
assign tree_c7       = {tree_s3 [64:0] & tree_s4 [64:0] | tree_s3 [64:0] & tree_s5 [64:0] | tree_s4 [64:0] & tree_s5 [64:0],1'b0};
assign tree_c8       = {tree_c0 [64:0] & tree_c1 [64:0] | tree_c0 [64:0] & tree_c2 [64:0] | tree_c1 [64:0] & tree_c2 [64:0],1'b0};
assign tree_c9       = {tree_c3 [64:0] & tree_c4 [64:0] | tree_c3 [64:0] & tree_c5 [64:0] | tree_c4 [64:0] & tree_c5 [64:0],1'b0};
assign tree_s0       = z0      & ~z1      & ~z2       | ~z0      & z1      & ~z2       | ~z0      & ~z1      & z2       | z0      & z1      & z2      ;
assign tree_s1       = z3      & ~z4      & ~z5       | ~z3      & z4      & ~z5       | ~z3      & ~z4      & z5       | z3      & z4      & z5      ;
assign tree_s10      = tree_s6 & ~tree_s7 & ~tree_s8  | ~tree_s6 & tree_s7 & ~tree_s8  | ~tree_s6 & ~tree_s7 & tree_s8  | tree_s6 & tree_s7 & tree_s8 ;
assign tree_s11      = tree_s9 & ~tree_c6 & ~tree_c7  | ~tree_s9 & tree_c6 & ~tree_c7  | ~tree_s9 & ~tree_c6 & tree_c7  | tree_s9 & tree_c6 & tree_c7 ;
assign tree_s12      = tree_c8 & ~tree_c9 & ~tree_s10 | ~tree_c8 & tree_c9 & ~tree_s10 | ~tree_c8 & ~tree_c9 & tree_s10 | tree_c8 & tree_c9 & tree_s10;
assign tree_s13      =  tree_s11 & ~tree_c10 & ~tree_c11
                     | ~tree_s11 &  tree_c10 & ~tree_c11
                     | ~tree_s11 & ~tree_c10 &  tree_c11
                     |  tree_s11 &  tree_c10 &  tree_c11;
assign tree_s14 =  tree_s12 & ~tree_s13 & ~tree_c12
                | ~tree_s12 &  tree_s13 & ~tree_c12
                | ~tree_s12 & ~tree_s13 &  tree_c12
                |  tree_s12 &  tree_s13 &  tree_c12;
assign tree_s15 =  tree_c13 & ~tree_s14 & ~tree_c14
                | ~tree_c13 &  tree_s14 & ~tree_c14
                | ~tree_c13 & ~tree_s14 &  tree_c14
                |  tree_c13 &  tree_s14 &  tree_c14;
assign tree_s2        = z6      & ~z7      & ~z8      | ~z6      & z7      & ~z8      | ~z6      & ~z7      & z8      | z6      & z7      & z8     ;
assign tree_s3        = z9      & ~z10     & ~z11     | ~z9      & z10     & ~z11     | ~z9      & ~z10     & z11     | z9      & z10     & z11    ;
assign tree_s4        = z12     & ~z13     & ~z14     | ~z12     & z13     & ~z14     | ~z12     & ~z13     & z14     | z12     & z13     & z14    ;
assign tree_s5        = z15     & ~z16     & ~z17     | ~z15     & z16     & ~z17     | ~z15     & ~z16     & z17     | z15     & z16     & z17    ;
assign tree_s6        = tree_s0 & ~tree_s1 & ~tree_s2 | ~tree_s0 & tree_s1 & ~tree_s2 | ~tree_s0 & ~tree_s1 & tree_s2 | tree_s0 & tree_s1 & tree_s2;
assign tree_s7        = tree_s3 & ~tree_s4 & ~tree_s5 | ~tree_s3 & tree_s4 & ~tree_s5 | ~tree_s3 & ~tree_s4 & tree_s5 | tree_s3 & tree_s4 & tree_s5;
assign tree_s8        = tree_c0 & ~tree_c1 & ~tree_c2 | ~tree_c0 & tree_c1 & ~tree_c2 | ~tree_c0 & ~tree_c1 & tree_c2 | tree_c0 & tree_c1 & tree_c2;
assign tree_s9        = tree_c3 & ~tree_c4 & ~tree_c5 | ~tree_c3 & tree_c4 & ~tree_c5 | ~tree_c3 & ~tree_c4 & tree_c5 | tree_c3 & tree_c4 & tree_c5;
assign u              = tree_c15;
assign v              = tree_s15;
assign y0             = {33{enc_neg[0 ]}} ^ b;
assign y1             = {33{enc_neg[1 ]}} ^ b;
assign y10            = {33{enc_neg[10]}} ^ b;
assign y11            = {33{enc_neg[11]}} ^ b;
assign y12            = {33{enc_neg[12]}} ^ b;
assign y13            = {33{enc_neg[13]}} ^ b;
assign y14            = {33{enc_neg[14]}} ^ b;
assign y15            = {33{enc_neg[15]}} ^ b;
assign y16            = {33{enc_neg[16]}} ^ b;
assign y2             = {33{enc_neg[2 ]}} ^ b;
assign y3             = {33{enc_neg[3 ]}} ^ b;
assign y4             = {33{enc_neg[4 ]}} ^ b;
assign y5             = {33{enc_neg[5 ]}} ^ b;
assign y6             = {33{enc_neg[6 ]}} ^ b;
assign y7             = {33{enc_neg[7 ]}} ^ b;
assign y8             = {33{enc_neg[8 ]}} ^ b;
assign y9             = {33{enc_neg[9 ]}} ^ b;
assign z0     [33:0 ] = {34{enc_m1[0]}} & {enc_lastb ^ enc_neg[0],y0} | {34{enc_m2[0]}} & {y0,enc_neg[0]};
assign z0     [65:34] = 32'h00000003;
assign z1     [35:2 ] = {34{enc_m1[1]}} & {enc_lastb ^ enc_neg[1],y1} | {34{enc_m2[1]}} & {y1,enc_neg[1]};
assign z1     [1 :0 ] = 2'h0        ;
assign z1     [65:36] = 30'h00000002;
assign z10    [53:20] = {34{enc_m1[10]}} & {enc_lastb ^ enc_neg[10],y10} | {34{enc_m2[10]}} & {y10,enc_neg[10]};
assign z10    [19:0 ] = 20'h00000;
assign z10    [65:54] = 12'h002  ;
assign z11    [55:22] = {34{enc_m1[11]}} & {enc_lastb ^ enc_neg[11],y11} | {34{enc_m2[11]}} & {y11,enc_neg[11]};
assign z11    [21:0 ] = 22'h000000;
assign z11    [65:56] = 10'h002   ;
assign z12    [57:24] = {34{enc_m1[12]}} & {enc_lastb ^ enc_neg[12],y12} | {34{enc_m2[12]}} & {y12,enc_neg[12]};
assign z12    [23:0 ] = 24'h000000;
assign z12    [65:58] = 8'h02     ;
assign z13    [59:26] = {34{enc_m1[13]}} & {enc_lastb ^ enc_neg[13],y13} | {34{enc_m2[13]}} & {y13,enc_neg[13]};
assign z13    [25:0 ] = 26'h0000000;
assign z13    [65:60] = 6'h02      ;
assign z14    [61:28] = {34{enc_m1[14]}} & {enc_lastb ^ enc_neg[14],y14} | {34{enc_m2[14]}} & {y14,enc_neg[14]};
assign z14    [27:0 ] = 28'h0000000;
assign z14    [65:62] = 4'h2       ;
assign z15    [63:30] = {34{enc_m1[15]}} & {enc_lastb ^ enc_neg[15],y15} | {34{enc_m2[15]}} & {y15,enc_neg[15]};
assign z15    [29:0 ] = 30'h00000000;
assign z15    [65:64] = 2'h2        ;
assign z16    [65:32] = {34{enc_m1[16]}} & {enc_lastb ^ enc_neg[16],y16} | {34{enc_m2[16]}} & {y16,enc_neg[16]};
assign z16    [31:0 ] = 32'h00000000;
assign z17    [   0 ] = enc_neg[0];
assign z17    [   1 ] = 1'h0;
assign z17    [   2 ] = enc_neg[1];
assign z17    [   3 ] = 1'h0;
assign z17    [   4 ] = enc_neg[2];
assign z17    [   5 ] = 1'h0;
assign z17    [   6 ] = enc_neg[3];
assign z17    [   7 ] = 1'h0;
assign z17    [   8 ] = enc_neg[4];
assign z17    [   9 ] = 1'h0;
assign z17    [   10] = enc_neg[5];
assign z17    [   11] = 1'h0;
assign z17    [   12] = enc_neg[6];
assign z17    [   13] = 1'h0;
assign z17    [   14] = enc_neg[7];
assign z17    [   15] = 1'h0;
assign z17    [   16] = enc_neg[8];
assign z17    [   17] = 1'h0;
assign z17    [   18] = enc_neg[9];
assign z17    [   19] = 1'h0;
assign z17    [   20] = enc_neg[10];
assign z17    [   21] = 1'h0;
assign z17    [   22] = enc_neg[11];
assign z17    [   23] = 1'h0;
assign z17    [   24] = enc_neg[12];
assign z17    [   25] = 1'h0;
assign z17    [   26] = enc_neg[13];
assign z17    [   27] = 1'h0;
assign z17    [   28] = enc_neg[14];
assign z17    [   29] = 1'h0;
assign z17    [   30] = enc_neg[15];
assign z17    [   31] = 1'h0;
assign z17    [   32] = enc_neg[16];
assign z17    [   33] = 1'h0;
assign z17    [   34] = !enc_ext[0];
assign z17    [   35] = 1'h0;
assign z17    [   36] = !enc_ext[1];
assign z17    [   37] = 1'h0;
assign z17    [   38] = !enc_ext[2];
assign z17    [   39] = 1'h0;
assign z17    [   40] = !enc_ext[3];
assign z17    [   41] = 1'h0;
assign z17    [   42] = !enc_ext[4];
assign z17    [   43] = 1'h0;
assign z17    [   44] = !enc_ext[5];
assign z17    [   45] = 1'h0;
assign z17    [   46] = !enc_ext[6];
assign z17    [   47] = 1'h0;
assign z17    [   48] = !enc_ext[7];
assign z17    [   49] = 1'h0;
assign z17    [   50] = !enc_ext[8];
assign z17    [   51] = 1'h0;
assign z17    [   52] = !enc_ext[9];
assign z17    [   53] = 1'h0;
assign z17    [   54] = !enc_ext[10];
assign z17    [   55] = 1'h0;
assign z17    [   56] = !enc_ext[11];
assign z17    [   57] = 1'h0;
assign z17    [   58] = !enc_ext[12];
assign z17    [   59] = 1'h0;
assign z17    [   60] = !enc_ext[13];
assign z17    [   61] = 1'h0;
assign z17    [   62] = !enc_ext[14];
assign z17    [   63] = 1'h0;
assign z17    [   64] = !enc_ext[15];
assign z17    [   65] = 1'h0;
assign z2     [37:4 ] = {34{enc_m1[2]}} & {enc_lastb ^ enc_neg[2],y2} | {34{enc_m2[2]}} & {y2,enc_neg[2]};
assign z2     [3 :0 ] = 4'h0       ;
assign z2     [65:38] = 28'h0000002;
assign z3     [39:6 ] = {34{enc_m1[3]}} & {enc_lastb ^ enc_neg[3],y3} | {34{enc_m2[3]}} & {y3,enc_neg[3]};
assign z3     [5 :0 ] = 6'h00      ;
assign z3     [65:40] = 26'h0000002;
assign z4     [41:8 ] = {34{enc_m1[4]}} & {enc_lastb ^ enc_neg[4],y4} | {34{enc_m2[4]}} & {y4,enc_neg[4]};
assign z4     [7 :0 ] = 8'h00     ;
assign z4     [65:42] = 24'h000002;
assign z5     [43:10] = {34{enc_m1[5]}} & {enc_lastb ^ enc_neg[5],y5} | {34{enc_m2[5]}} & {y5,enc_neg[5]};
assign z5     [9 :0 ] = 10'h000   ;
assign z5     [65:44] = 22'h000002;
assign z6     [45:12] = {34{enc_m1[6]}} & {enc_lastb ^ enc_neg[6],y6} | {34{enc_m2[6]}} & {y6,enc_neg[6]};
assign z6     [11:0 ] = 12'h000  ;
assign z6     [65:46] = 20'h00002;
assign z7     [47:14] = {34{enc_m1[7]}} & {enc_lastb ^ enc_neg[7],y7} | {34{enc_m2[7]}} & {y7,enc_neg[7]};
assign z7     [13:0 ] = 14'h0000 ;
assign z7     [65:48] = 18'h00002;
assign z8     [49:16] = {34{enc_m1[8]}} & {enc_lastb ^ enc_neg[8],y8} | {34{enc_m2[8]}} & {y8,enc_neg[8]};
assign z8     [15:0 ] = 16'h0000;
assign z8     [65:50] = 16'h0002;
assign z9     [51:18] = {34{enc_m1[9]}} & {enc_lastb ^ enc_neg[9],y9} | {34{enc_m2[9]}} & {y9,enc_neg[9]};
assign z9     [17:0 ] = 18'h00000;
assign z9     [65:52] = 14'h0002 ;

endmodule // mul
